module computer(input clk, reset, input[1023 : 0] code);

endmodule
